module dec2to4 ( 
	a,
	e,
	o
	) ;

input [1:0] a;
input  e;
inout [3:0] o;
