module entalu3bits ( 
	a,
	b,
	oper,
	result
	) ;

input [2:0] a;
input [2:0] b;
input [1:0] oper;
inout [3:0] result;
