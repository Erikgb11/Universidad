module ula ( 
	a,
	b,
	o,
	sel
	) ;

input [3:0] a;
input [3:0] b;
inout [3:0] o;
input [2:0] sel;
